`timescale 1ns / 1ps

module decoder(
    input [31:0] instruction,
    output [1:0] instr_type,
    output [2:0] data_instr_type
    );


endmodule
